VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM8
  CLASS BLOCK ;
  FOREIGN RAM8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 108.100 BY 21.760 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.100 5.480 108.100 6.080 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.100 8.200 108.100 8.800 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.100 10.920 108.100 11.520 ;
    END
  END A0[2]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.100 13.640 108.100 14.240 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.000 ;
    END
  END Di0[0]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 2.000 ;
    END
  END Di0[1]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.000 ;
    END
  END Di0[2]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.000 ;
    END
  END Di0[7]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 19.760 7.270 21.760 ;
    END
  END Do0[0]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 19.760 20.610 21.760 ;
    END
  END Do0[1]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 19.760 33.950 21.760 ;
    END
  END Do0[2]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 19.760 47.290 21.760 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 19.760 60.630 21.760 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 19.760 73.970 21.760 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 19.760 87.310 21.760 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 19.760 100.650 21.760 ;
    END
  END Do0[7]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.100 2.760 108.100 3.360 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.320 -0.240 93.920 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.145 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 -0.240 108.100 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 0.145 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 5.200 108.100 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 10.640 0.145 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 10.640 108.100 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 16.080 0.145 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 16.080 108.100 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 21.520 0.145 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 21.520 108.100 22.000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.520 -0.240 17.120 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.145 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 2.480 108.100 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 7.920 0.145 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 7.920 108.100 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 13.360 0.145 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 13.360 108.100 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 18.800 0.145 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 107.955 18.800 108.100 19.280 ;
    END
  END VPWR
  PIN WE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.100 16.360 108.100 16.960 ;
    END
  END WE0
  OBS
      LAYER pwell ;
        RECT 0.605 21.655 0.775 21.845 ;
        RECT 6.130 21.655 6.300 21.845 ;
        RECT 10.725 21.655 10.895 21.845 ;
        RECT 16.250 21.655 16.420 21.845 ;
        RECT 20.845 21.655 21.015 21.845 ;
        RECT 26.370 21.655 26.540 21.845 ;
        RECT 30.965 21.655 31.135 21.845 ;
        RECT 36.490 21.655 36.660 21.845 ;
        RECT 41.085 21.655 41.255 21.845 ;
        RECT 46.610 21.655 46.780 21.845 ;
        RECT 51.205 21.655 51.375 21.845 ;
        RECT 56.730 21.655 56.900 21.845 ;
        RECT 61.325 21.655 61.495 21.845 ;
        RECT 66.850 21.655 67.020 21.845 ;
        RECT 71.445 21.655 71.615 21.845 ;
        RECT 76.970 21.655 77.140 21.845 ;
        RECT 81.570 21.655 81.740 21.845 ;
        RECT 88.005 21.675 88.175 21.845 ;
        RECT 90.305 21.695 90.475 21.845 ;
        RECT 91.225 21.675 91.395 21.845 ;
        RECT 92.605 21.675 92.775 21.845 ;
        RECT 94.445 21.655 94.615 21.845 ;
        RECT 97.205 21.655 97.375 21.845 ;
        RECT 99.505 21.655 99.675 21.845 ;
        RECT 100.890 21.655 101.060 21.845 ;
        RECT 105.025 21.655 105.195 21.845 ;
      LAYER nwell ;
        RECT -0.190 20.405 82.415 20.455 ;
        RECT 84.040 20.405 108.290 20.455 ;
        RECT -0.190 17.675 108.290 20.405 ;
        RECT -0.190 17.625 81.955 17.675 ;
        RECT 83.580 17.625 108.290 17.675 ;
        RECT -0.190 14.965 82.415 15.015 ;
        RECT 84.040 14.965 108.290 15.015 ;
        RECT -0.190 12.235 108.290 14.965 ;
        RECT -0.190 12.185 81.955 12.235 ;
        RECT 83.580 12.185 108.290 12.235 ;
        RECT -0.190 9.525 82.415 9.575 ;
        RECT 84.040 9.525 108.290 9.575 ;
        RECT -0.190 6.795 108.290 9.525 ;
        RECT -0.190 6.745 81.955 6.795 ;
        RECT 83.580 6.745 108.290 6.795 ;
        RECT -0.190 4.085 82.415 4.135 ;
        RECT 84.040 4.085 108.290 4.135 ;
        RECT -0.190 1.355 108.290 4.085 ;
        RECT -0.190 1.305 81.955 1.355 ;
        RECT 83.580 1.305 108.290 1.355 ;
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 5.670 -0.085 5.840 0.105 ;
        RECT 10.265 -0.085 10.435 0.105 ;
        RECT 15.790 -0.085 15.960 0.105 ;
        RECT 20.385 -0.085 20.555 0.105 ;
        RECT 25.910 -0.085 26.080 0.105 ;
        RECT 30.505 -0.085 30.675 0.105 ;
        RECT 36.030 -0.085 36.200 0.105 ;
        RECT 40.625 -0.085 40.795 0.105 ;
        RECT 46.150 -0.085 46.320 0.105 ;
        RECT 50.745 -0.085 50.915 0.105 ;
        RECT 56.270 -0.085 56.440 0.105 ;
        RECT 60.865 -0.085 61.035 0.105 ;
        RECT 66.390 -0.085 66.560 0.105 ;
        RECT 70.985 -0.085 71.155 0.105 ;
        RECT 76.510 -0.085 76.680 0.105 ;
        RECT 81.110 -0.085 81.280 0.105 ;
        RECT 87.545 -0.085 87.715 0.085 ;
        RECT 89.845 -0.085 90.015 0.065 ;
        RECT 90.765 -0.085 90.935 0.085 ;
        RECT 92.145 -0.085 92.315 0.085 ;
        RECT 93.985 -0.085 94.155 0.105 ;
        RECT 96.745 -0.085 96.915 0.105 ;
        RECT 99.045 -0.085 99.215 0.105 ;
        RECT 100.885 -0.085 101.055 0.105 ;
        RECT 106.405 -0.085 106.575 0.105 ;
      LAYER li1 ;
        RECT 0.000 21.675 108.100 21.845 ;
      LAYER li1 ;
        RECT 0.000 0.085 108.100 21.675 ;
      LAYER li1 ;
        RECT 0.000 -0.085 108.100 0.085 ;
      LAYER met1 ;
        RECT 0.145 21.675 107.955 22.000 ;
        RECT 0.425 21.240 107.675 21.675 ;
        RECT 0.085 19.560 107.955 21.240 ;
        RECT 0.425 18.520 107.675 19.560 ;
        RECT 0.085 16.840 107.955 18.520 ;
        RECT 0.425 15.800 107.675 16.840 ;
        RECT 0.085 14.120 107.955 15.800 ;
        RECT 0.425 13.080 107.675 14.120 ;
        RECT 0.085 11.400 107.955 13.080 ;
        RECT 0.425 10.360 107.675 11.400 ;
        RECT 0.085 8.680 107.955 10.360 ;
        RECT 0.425 7.640 107.675 8.680 ;
        RECT 0.085 5.960 107.955 7.640 ;
        RECT 0.425 4.920 107.675 5.960 ;
        RECT 0.085 3.240 107.955 4.920 ;
        RECT 0.425 2.200 107.675 3.240 ;
        RECT 0.085 0.520 107.955 2.200 ;
        RECT 0.425 0.085 107.675 0.520 ;
        RECT 0.145 -0.240 107.955 0.085 ;
      LAYER met2 ;
        RECT 92.350 21.760 93.890 21.945 ;
        RECT 1.940 19.480 6.710 21.760 ;
        RECT 7.550 19.480 20.050 21.760 ;
        RECT 20.890 19.480 33.390 21.760 ;
        RECT 34.230 19.480 46.730 21.760 ;
        RECT 47.570 19.480 60.070 21.760 ;
        RECT 60.910 19.480 73.410 21.760 ;
        RECT 74.250 19.480 86.750 21.760 ;
        RECT 87.590 19.480 100.090 21.760 ;
        RECT 100.930 19.480 106.160 21.760 ;
        RECT 1.940 2.280 106.160 19.480 ;
        RECT 1.940 0.000 6.710 2.280 ;
        RECT 7.550 0.000 20.050 2.280 ;
        RECT 20.890 0.000 33.390 2.280 ;
        RECT 34.230 0.000 46.730 2.280 ;
        RECT 47.570 0.000 60.070 2.280 ;
        RECT 60.910 0.000 73.410 2.280 ;
        RECT 74.250 0.000 86.750 2.280 ;
        RECT 87.590 0.000 100.090 2.280 ;
        RECT 100.930 0.000 106.160 2.280 ;
        RECT 92.350 -0.185 93.890 0.000 ;
      LAYER met3 ;
        RECT 92.330 21.760 93.910 21.925 ;
        RECT 15.530 17.360 106.100 21.760 ;
        RECT 15.530 15.960 105.700 17.360 ;
        RECT 15.530 14.640 106.100 15.960 ;
        RECT 15.530 13.240 105.700 14.640 ;
        RECT 15.530 11.920 106.100 13.240 ;
        RECT 15.530 10.520 105.700 11.920 ;
        RECT 15.530 9.200 106.100 10.520 ;
        RECT 15.530 7.800 105.700 9.200 ;
        RECT 15.530 6.480 106.100 7.800 ;
        RECT 15.530 5.080 105.700 6.480 ;
        RECT 15.530 3.760 106.100 5.080 ;
        RECT 15.530 2.360 105.700 3.760 ;
        RECT 15.530 0.000 106.100 2.360 ;
        RECT 92.330 -0.165 93.910 0.000 ;
  END
END RAM8
END LIBRARY

