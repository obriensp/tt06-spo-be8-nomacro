VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO I2C
  CLASS BLOCK ;
  FOREIGN I2C ;
  ORIGIN -2.760 0.000 ;
  SIZE 155.480 BY 32.640 ;
  PIN PADDR[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 132.790 0.000 133.090 1.000 ;
    END
  END PADDR[0]
  PIN PADDR[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 129.110 0.000 129.410 4.570 ;
    END
  END PADDR[1]
  PIN PADDR[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 125.430 0.000 125.730 1.000 ;
    END
  END PADDR[2]
  PIN PADDR[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 121.750 0.000 122.050 3.890 ;
    END
  END PADDR[3]
  PIN PADDR[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 118.070 0.000 118.370 1.000 ;
    END
  END PADDR[4]
  PIN PCLK
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 154.870 0.000 155.170 1.000 ;
    END
  END PCLK
  PIN PENABLE
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 103.350 0.000 103.650 1.000 ;
    END
  END PENABLE
  PIN PRDATA[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 48.150 0.000 48.450 5.930 ;
    END
  END PRDATA[0]
  PIN PRDATA[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 44.470 0.000 44.770 4.960 ;
    END
  END PRDATA[1]
  PIN PRDATA[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 40.790 0.000 41.090 1.000 ;
    END
  END PRDATA[2]
  PIN PRDATA[3]
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 37.110 0.000 37.410 1.000 ;
    END
  END PRDATA[3]
  PIN PRDATA[4]
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 33.430 0.000 33.730 1.000 ;
    END
  END PRDATA[4]
  PIN PRDATA[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 29.750 0.000 30.050 1.000 ;
    END
  END PRDATA[5]
  PIN PRDATA[6]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 26.070 0.000 26.370 1.000 ;
    END
  END PRDATA[6]
  PIN PRDATA[7]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 22.390 0.000 22.690 4.570 ;
    END
  END PRDATA[7]
  PIN PREADY
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 3.990 0.000 4.290 1.000 ;
    END
  END PREADY
  PIN PRESETn
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 151.190 0.000 151.490 1.000 ;
    END
  END PRESETn
  PIN PSEL
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 147.510 0.000 147.810 1.000 ;
    END
  END PSEL
  PIN PWDATA[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.950 0.000 85.250 1.000 ;
    END
  END PWDATA[0]
  PIN PWDATA[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 81.270 0.000 81.570 1.000 ;
    END
  END PWDATA[1]
  PIN PWDATA[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 77.590 0.000 77.890 1.000 ;
    END
  END PWDATA[2]
  PIN PWDATA[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 73.910 0.000 74.210 1.000 ;
    END
  END PWDATA[3]
  PIN PWDATA[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 70.230 0.000 70.530 1.000 ;
    END
  END PWDATA[4]
  PIN PWDATA[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 66.550 0.000 66.850 3.890 ;
    END
  END PWDATA[5]
  PIN PWDATA[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 62.870 0.000 63.170 1.000 ;
    END
  END PWDATA[6]
  PIN PWDATA[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 59.190 0.000 59.490 1.000 ;
    END
  END PWDATA[7]
  PIN PWRITE
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 99.670 0.000 99.970 1.000 ;
    END
  END PWRITE
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2.760 29.680 2.905 30.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 30.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 2.480 2.905 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 2.480 158.240 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 7.920 2.905 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 7.920 158.240 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 13.360 2.905 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 13.360 158.240 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 18.800 2.905 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 18.800 158.240 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 24.240 2.905 24.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 24.240 158.240 24.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 29.680 158.240 30.160 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 158.095 16.080 158.240 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 26.960 158.240 27.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 26.960 2.905 27.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 21.520 158.240 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 21.520 2.905 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 16.080 2.905 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 10.640 158.240 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 10.640 2.905 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 158.095 5.200 158.240 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.760 5.200 2.905 5.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 30.160 ;
    END
  END VPWR
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 153.870 28.750 154.170 32.640 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met3 ;
        RECT 157.550 31.640 157.850 32.640 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 150.190 31.640 150.490 32.640 ;
    END
  END rst_n
  PIN ui_in[0]
    PORT
      LAYER met3 ;
        RECT 146.510 31.640 146.810 32.640 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met3 ;
        RECT 142.830 31.640 143.130 32.640 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met3 ;
        RECT 139.150 31.640 139.450 32.640 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met3 ;
        RECT 135.470 31.640 135.770 32.640 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met3 ;
        RECT 131.790 31.640 132.090 32.640 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met3 ;
        RECT 128.110 31.640 128.410 32.640 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met3 ;
        RECT 124.430 31.640 124.730 32.640 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met3 ;
        RECT 120.750 31.640 121.050 32.640 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met3 ;
        RECT 117.070 31.640 117.370 32.640 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met3 ;
        RECT 113.390 31.640 113.690 32.640 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 109.710 30.110 110.010 32.640 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 106.030 31.640 106.330 32.640 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met3 ;
        RECT 102.350 31.640 102.650 32.640 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met3 ;
        RECT 98.670 31.640 98.970 32.640 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met3 ;
        RECT 94.990 31.640 95.290 32.640 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met3 ;
        RECT 91.310 31.640 91.610 32.640 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 28.750 31.640 29.050 32.640 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 25.070 31.640 25.370 32.640 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 21.390 31.640 21.690 32.640 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 17.710 31.640 18.010 32.640 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 14.030 31.640 14.330 32.640 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 10.350 31.640 10.650 32.640 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 6.670 31.640 6.970 32.640 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2.990 31.640 3.290 32.640 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.190 31.640 58.490 32.640 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 54.510 31.640 54.810 32.640 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 50.830 31.640 51.130 32.640 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 47.150 31.640 47.450 32.640 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 43.470 31.640 43.770 32.640 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 39.790 31.640 40.090 32.640 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 36.110 31.640 36.410 32.640 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 32.430 31.640 32.730 32.640 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 87.630 31.640 87.930 32.640 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 83.950 31.640 84.250 32.640 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 80.270 31.640 80.570 32.640 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.590 31.640 76.890 32.640 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 72.910 31.640 73.210 32.640 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 69.230 31.640 69.530 32.640 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 65.550 31.640 65.850 32.640 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 61.870 31.640 62.170 32.640 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 25.785 158.430 28.615 ;
        RECT 2.570 20.345 158.430 23.175 ;
        RECT 2.570 14.905 158.430 17.735 ;
        RECT 2.570 9.465 158.430 12.295 ;
        RECT 2.570 4.025 158.430 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 158.240 30.005 ;
      LAYER met1 ;
        RECT 2.905 30.440 158.095 31.240 ;
        RECT 3.185 29.400 157.815 30.440 ;
        RECT 2.905 27.720 158.095 29.400 ;
        RECT 3.185 26.680 157.815 27.720 ;
        RECT 2.905 25.000 158.095 26.680 ;
        RECT 3.185 23.960 157.815 25.000 ;
        RECT 2.905 22.280 158.095 23.960 ;
        RECT 3.185 21.240 157.815 22.280 ;
        RECT 2.905 19.560 158.095 21.240 ;
        RECT 3.185 18.520 157.815 19.560 ;
        RECT 2.905 16.840 158.095 18.520 ;
        RECT 3.185 15.800 157.815 16.840 ;
        RECT 2.905 14.120 158.095 15.800 ;
        RECT 3.185 13.080 157.815 14.120 ;
        RECT 2.905 11.400 158.095 13.080 ;
        RECT 3.185 10.360 157.815 11.400 ;
        RECT 2.905 8.680 158.095 10.360 ;
        RECT 3.185 7.640 157.815 8.680 ;
        RECT 2.905 5.960 158.095 7.640 ;
        RECT 3.185 4.920 157.815 5.960 ;
        RECT 2.905 3.240 158.095 4.920 ;
        RECT 3.185 2.200 157.815 3.240 ;
        RECT 2.905 0.380 158.095 2.200 ;
      LAYER met2 ;
        RECT 4.690 0.155 156.300 32.485 ;
      LAYER met3 ;
        RECT 3.690 31.240 6.270 32.465 ;
        RECT 7.370 31.240 9.950 32.465 ;
        RECT 11.050 31.240 13.630 32.465 ;
        RECT 14.730 31.240 17.310 32.465 ;
        RECT 18.410 31.240 20.990 32.465 ;
        RECT 22.090 31.240 24.670 32.465 ;
        RECT 25.770 31.240 28.350 32.465 ;
        RECT 29.450 31.240 32.030 32.465 ;
        RECT 33.130 31.240 35.710 32.465 ;
        RECT 36.810 31.240 39.390 32.465 ;
        RECT 40.490 31.240 43.070 32.465 ;
        RECT 44.170 31.240 46.750 32.465 ;
        RECT 47.850 31.240 50.430 32.465 ;
        RECT 51.530 31.240 54.110 32.465 ;
        RECT 55.210 31.240 57.790 32.465 ;
        RECT 58.890 31.240 61.470 32.465 ;
        RECT 62.570 31.240 65.150 32.465 ;
        RECT 66.250 31.240 68.830 32.465 ;
        RECT 69.930 31.240 72.510 32.465 ;
        RECT 73.610 31.240 76.190 32.465 ;
        RECT 77.290 31.240 79.870 32.465 ;
        RECT 80.970 31.240 83.550 32.465 ;
        RECT 84.650 31.240 87.230 32.465 ;
        RECT 88.330 31.240 90.910 32.465 ;
        RECT 92.010 31.240 94.590 32.465 ;
        RECT 95.690 31.240 98.270 32.465 ;
        RECT 99.370 31.240 101.950 32.465 ;
        RECT 103.050 31.240 105.630 32.465 ;
        RECT 106.730 31.240 109.310 32.465 ;
        RECT 3.290 29.710 109.310 31.240 ;
        RECT 110.410 31.240 112.990 32.465 ;
        RECT 114.090 31.240 116.670 32.465 ;
        RECT 117.770 31.240 120.350 32.465 ;
        RECT 121.450 31.240 124.030 32.465 ;
        RECT 125.130 31.240 127.710 32.465 ;
        RECT 128.810 31.240 131.390 32.465 ;
        RECT 132.490 31.240 135.070 32.465 ;
        RECT 136.170 31.240 138.750 32.465 ;
        RECT 139.850 31.240 142.430 32.465 ;
        RECT 143.530 31.240 146.110 32.465 ;
        RECT 147.210 31.240 149.790 32.465 ;
        RECT 150.890 31.240 153.470 32.465 ;
        RECT 110.410 29.710 153.470 31.240 ;
        RECT 3.290 28.350 153.470 29.710 ;
        RECT 154.570 28.350 155.875 32.465 ;
        RECT 3.290 6.330 155.875 28.350 ;
        RECT 3.290 5.360 47.750 6.330 ;
        RECT 3.290 4.970 44.070 5.360 ;
        RECT 3.290 1.400 21.990 4.970 ;
        RECT 3.290 0.175 3.590 1.400 ;
        RECT 4.690 0.175 21.990 1.400 ;
        RECT 23.090 1.400 44.070 4.970 ;
        RECT 23.090 0.175 25.670 1.400 ;
        RECT 26.770 0.175 29.350 1.400 ;
        RECT 30.450 0.175 33.030 1.400 ;
        RECT 34.130 0.175 36.710 1.400 ;
        RECT 37.810 0.175 40.390 1.400 ;
        RECT 41.490 0.175 44.070 1.400 ;
        RECT 45.170 0.175 47.750 5.360 ;
        RECT 48.850 4.970 155.875 6.330 ;
        RECT 48.850 4.290 128.710 4.970 ;
        RECT 48.850 1.400 66.150 4.290 ;
        RECT 48.850 0.175 58.790 1.400 ;
        RECT 59.890 0.175 62.470 1.400 ;
        RECT 63.570 0.175 66.150 1.400 ;
        RECT 67.250 1.400 121.350 4.290 ;
        RECT 67.250 0.175 69.830 1.400 ;
        RECT 70.930 0.175 73.510 1.400 ;
        RECT 74.610 0.175 77.190 1.400 ;
        RECT 78.290 0.175 80.870 1.400 ;
        RECT 81.970 0.175 84.550 1.400 ;
        RECT 85.650 0.175 99.270 1.400 ;
        RECT 100.370 0.175 102.950 1.400 ;
        RECT 104.050 0.175 117.670 1.400 ;
        RECT 118.770 0.175 121.350 1.400 ;
        RECT 122.450 1.400 128.710 4.290 ;
        RECT 122.450 0.175 125.030 1.400 ;
        RECT 126.130 0.175 128.710 1.400 ;
        RECT 129.810 1.400 155.875 4.970 ;
        RECT 129.810 0.175 132.390 1.400 ;
        RECT 133.490 0.175 147.110 1.400 ;
        RECT 148.210 0.175 150.790 1.400 ;
        RECT 151.890 0.175 154.470 1.400 ;
        RECT 155.570 0.175 155.875 1.400 ;
      LAYER met4 ;
        RECT 73.895 7.655 86.185 19.545 ;
  END
END I2C
END LIBRARY

