VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM8
  CLASS BLOCK ;
  FOREIGN RAM8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 121.440 BY 21.760 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.440 5.480 121.440 6.080 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.440 8.200 121.440 8.800 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.440 10.920 121.440 11.520 ;
    END
  END A0[2]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.440 13.640 121.440 14.240 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.000 ;
    END
  END Di0[0]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.000 ;
    END
  END Di0[1]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 2.000 ;
    END
  END Di0[2]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.000 ;
    END
  END Di0[7]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 19.760 7.730 21.760 ;
    END
  END Do0[0]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 19.760 22.910 21.760 ;
    END
  END Do0[1]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 19.760 38.090 21.760 ;
    END
  END Do0[2]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 19.760 53.270 21.760 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 19.760 68.450 21.760 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 19.760 83.630 21.760 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 19.760 98.810 21.760 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 19.760 113.990 21.760 ;
    END
  END Do0[7]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.440 2.760 121.440 3.360 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.320 -0.240 93.920 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.145 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 -0.240 121.440 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 0.145 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 5.200 121.440 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 10.640 0.145 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 10.640 121.440 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 16.080 0.145 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 16.080 121.440 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 21.520 0.145 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 21.520 121.440 22.000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.520 -0.240 17.120 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.145 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 2.480 121.440 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 7.920 0.145 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 7.920 121.440 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 13.360 0.145 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 13.360 121.440 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 18.800 0.145 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 121.295 18.800 121.440 19.280 ;
    END
  END VPWR
  PIN WE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.440 16.360 121.440 16.960 ;
    END
  END WE0
  OBS
      LAYER pwell ;
        RECT 0.605 21.655 0.775 21.845 ;
        RECT 7.970 21.655 8.140 21.845 ;
        RECT 12.565 21.655 12.735 21.845 ;
        RECT 19.930 21.655 20.100 21.845 ;
        RECT 24.525 21.655 24.695 21.845 ;
        RECT 31.890 21.655 32.060 21.845 ;
        RECT 36.485 21.655 36.655 21.845 ;
        RECT 43.850 21.655 44.020 21.845 ;
        RECT 48.445 21.655 48.615 21.845 ;
        RECT 55.810 21.655 55.980 21.845 ;
        RECT 60.405 21.655 60.575 21.845 ;
        RECT 67.770 21.655 67.940 21.845 ;
        RECT 72.365 21.655 72.535 21.845 ;
        RECT 79.730 21.655 79.900 21.845 ;
        RECT 84.325 21.655 84.495 21.845 ;
        RECT 91.690 21.655 91.860 21.845 ;
        RECT 96.290 21.655 96.460 21.845 ;
        RECT 102.725 21.675 102.895 21.845 ;
        RECT 105.025 21.695 105.195 21.845 ;
        RECT 105.945 21.675 106.115 21.845 ;
        RECT 107.325 21.655 107.495 21.845 ;
        RECT 110.545 21.655 110.715 21.845 ;
        RECT 112.845 21.655 113.015 21.845 ;
        RECT 114.230 21.655 114.400 21.845 ;
        RECT 118.365 21.655 118.535 21.845 ;
      LAYER nwell ;
        RECT -0.190 20.405 97.135 20.455 ;
        RECT 98.760 20.405 121.630 20.455 ;
        RECT -0.190 17.675 121.630 20.405 ;
        RECT -0.190 17.625 96.675 17.675 ;
        RECT 98.300 17.625 121.630 17.675 ;
        RECT -0.190 14.965 97.135 15.015 ;
        RECT 98.760 14.965 121.630 15.015 ;
        RECT -0.190 12.235 121.630 14.965 ;
        RECT -0.190 12.185 96.675 12.235 ;
        RECT 98.300 12.185 121.630 12.235 ;
        RECT -0.190 9.525 97.135 9.575 ;
        RECT 98.760 9.525 121.630 9.575 ;
        RECT -0.190 6.795 121.630 9.525 ;
        RECT -0.190 6.745 96.675 6.795 ;
        RECT 98.300 6.745 121.630 6.795 ;
        RECT -0.190 4.085 97.135 4.135 ;
        RECT 98.760 4.085 121.630 4.135 ;
        RECT -0.190 1.355 121.630 4.085 ;
        RECT -0.190 1.305 96.675 1.355 ;
        RECT 98.300 1.305 121.630 1.355 ;
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 7.510 -0.085 7.680 0.105 ;
        RECT 12.105 -0.085 12.275 0.105 ;
        RECT 19.470 -0.085 19.640 0.105 ;
        RECT 24.065 -0.085 24.235 0.105 ;
        RECT 31.430 -0.085 31.600 0.105 ;
        RECT 36.025 -0.085 36.195 0.105 ;
        RECT 43.390 -0.085 43.560 0.105 ;
        RECT 47.985 -0.085 48.155 0.105 ;
        RECT 55.350 -0.085 55.520 0.105 ;
        RECT 59.945 -0.085 60.115 0.105 ;
        RECT 67.310 -0.085 67.480 0.105 ;
        RECT 71.905 -0.085 72.075 0.105 ;
        RECT 79.270 -0.085 79.440 0.105 ;
        RECT 83.865 -0.085 84.035 0.105 ;
        RECT 91.230 -0.085 91.400 0.105 ;
        RECT 95.830 -0.085 96.000 0.105 ;
        RECT 102.265 -0.085 102.435 0.085 ;
        RECT 104.565 -0.085 104.735 0.065 ;
        RECT 105.485 -0.085 105.655 0.085 ;
        RECT 106.865 -0.085 107.035 0.105 ;
        RECT 110.085 -0.085 110.255 0.105 ;
        RECT 112.385 -0.085 112.555 0.105 ;
        RECT 114.225 -0.085 114.395 0.105 ;
        RECT 119.745 -0.085 119.915 0.105 ;
      LAYER li1 ;
        RECT 0.000 21.675 121.440 21.845 ;
      LAYER li1 ;
        RECT 0.000 0.085 121.440 21.675 ;
      LAYER li1 ;
        RECT 0.000 -0.085 121.440 0.085 ;
      LAYER met1 ;
        RECT 0.145 21.675 121.295 22.000 ;
        RECT 0.425 21.240 121.015 21.675 ;
        RECT 0.085 19.560 121.295 21.240 ;
        RECT 0.425 18.520 121.015 19.560 ;
        RECT 0.085 16.840 121.295 18.520 ;
        RECT 0.425 15.800 121.015 16.840 ;
        RECT 0.085 14.120 121.295 15.800 ;
        RECT 0.425 13.080 121.015 14.120 ;
        RECT 0.085 11.400 121.295 13.080 ;
        RECT 0.425 10.360 121.015 11.400 ;
        RECT 0.085 8.680 121.295 10.360 ;
        RECT 0.425 7.640 121.015 8.680 ;
        RECT 0.085 5.960 121.295 7.640 ;
        RECT 0.425 4.920 121.015 5.960 ;
        RECT 0.085 3.240 121.295 4.920 ;
        RECT 0.425 2.200 121.015 3.240 ;
        RECT 0.085 0.520 121.295 2.200 ;
        RECT 0.425 0.085 121.015 0.520 ;
        RECT 0.145 -0.240 121.295 0.085 ;
      LAYER met2 ;
        RECT 92.350 21.760 93.890 21.945 ;
        RECT 1.940 19.480 7.170 21.760 ;
        RECT 8.010 19.480 22.350 21.760 ;
        RECT 23.190 19.480 37.530 21.760 ;
        RECT 38.370 19.480 52.710 21.760 ;
        RECT 53.550 19.480 67.890 21.760 ;
        RECT 68.730 19.480 83.070 21.760 ;
        RECT 83.910 19.480 98.250 21.760 ;
        RECT 99.090 19.480 113.430 21.760 ;
        RECT 114.270 19.480 119.050 21.760 ;
        RECT 1.940 2.280 119.050 19.480 ;
        RECT 1.940 0.000 7.170 2.280 ;
        RECT 8.010 0.000 22.350 2.280 ;
        RECT 23.190 0.000 37.530 2.280 ;
        RECT 38.370 0.000 52.710 2.280 ;
        RECT 53.550 0.000 67.890 2.280 ;
        RECT 68.730 0.000 83.070 2.280 ;
        RECT 83.910 0.000 98.250 2.280 ;
        RECT 99.090 0.000 113.430 2.280 ;
        RECT 114.270 0.000 119.050 2.280 ;
        RECT 92.350 -0.185 93.890 0.000 ;
      LAYER met3 ;
        RECT 92.330 21.760 93.910 21.925 ;
        RECT 15.530 17.360 119.440 21.760 ;
        RECT 15.530 15.960 119.040 17.360 ;
        RECT 15.530 14.640 119.440 15.960 ;
        RECT 15.530 13.240 119.040 14.640 ;
        RECT 15.530 11.920 119.440 13.240 ;
        RECT 15.530 10.520 119.040 11.920 ;
        RECT 15.530 9.200 119.440 10.520 ;
        RECT 15.530 7.800 119.040 9.200 ;
        RECT 15.530 6.480 119.440 7.800 ;
        RECT 15.530 5.080 119.040 6.480 ;
        RECT 15.530 3.760 119.440 5.080 ;
        RECT 15.530 2.360 119.040 3.760 ;
        RECT 15.530 0.000 119.440 2.360 ;
        RECT 92.330 -0.165 93.910 0.000 ;
  END
END RAM8
END LIBRARY

