VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM16
  CLASS BLOCK ;
  FOREIGN RAM16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 124.660 BY 43.520 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.660 9.560 124.660 10.160 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.660 15.000 124.660 15.600 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.660 20.440 124.660 21.040 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.660 25.880 124.660 26.480 ;
    END
  END A0[3]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.660 31.320 124.660 31.920 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 41.520 7.270 43.520 ;
    END
  END Di0[0]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 41.520 14.630 43.520 ;
    END
  END Di0[1]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 41.520 21.990 43.520 ;
    END
  END Di0[2]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 41.520 29.350 43.520 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 41.520 36.710 43.520 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 41.520 44.070 43.520 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 41.520 51.430 43.520 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 41.520 58.790 43.520 ;
    END
  END Di0[7]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 41.520 66.150 43.520 ;
    END
  END Do0[0]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 41.520 73.510 43.520 ;
    END
  END Do0[1]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 41.520 80.870 43.520 ;
    END
  END Do0[2]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 41.520 88.230 43.520 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 41.520 95.590 43.520 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 41.520 102.950 43.520 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 41.520 110.310 43.520 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 41.520 117.670 43.520 ;
    END
  END Do0[7]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.660 4.120 124.660 4.720 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.120 -0.240 42.720 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.320 -0.240 93.920 43.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.145 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 -0.240 124.660 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 0.145 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 5.200 124.660 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 10.640 0.145 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 10.640 124.660 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 16.080 0.145 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 16.080 124.660 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 21.520 0.145 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 21.520 124.660 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 26.960 0.145 27.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 26.960 124.660 27.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 32.400 0.145 32.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 32.400 124.660 32.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 37.840 0.145 38.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 37.840 124.660 38.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 43.280 0.145 43.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 43.280 124.660 43.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.520 -0.240 17.120 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.720 -0.240 68.320 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.920 -0.240 119.520 43.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.145 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 2.480 124.660 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 7.920 0.145 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 7.920 124.660 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 13.360 0.145 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 13.360 124.660 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 18.800 0.145 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 18.800 124.660 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 24.240 0.145 24.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 24.240 124.660 24.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 29.680 0.145 30.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 29.680 124.660 30.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 35.120 0.145 35.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 35.120 124.660 35.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 40.560 0.145 41.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 124.515 40.560 124.660 41.040 ;
    END
  END VPWR
  PIN WE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.660 36.760 124.660 37.360 ;
    END
  END WE0
  OBS
      LAYER pwell ;
        RECT 0.605 43.415 0.775 43.605 ;
        RECT 7.970 43.415 8.140 43.605 ;
        RECT 12.565 43.415 12.735 43.605 ;
        RECT 19.930 43.415 20.100 43.605 ;
        RECT 24.525 43.415 24.695 43.605 ;
        RECT 31.890 43.415 32.060 43.605 ;
        RECT 36.485 43.415 36.655 43.605 ;
        RECT 43.850 43.415 44.020 43.605 ;
        RECT 48.445 43.415 48.615 43.605 ;
        RECT 55.810 43.415 55.980 43.605 ;
        RECT 60.405 43.415 60.575 43.605 ;
        RECT 67.770 43.415 67.940 43.605 ;
        RECT 72.365 43.415 72.535 43.605 ;
        RECT 79.730 43.415 79.900 43.605 ;
        RECT 84.325 43.415 84.495 43.605 ;
        RECT 91.690 43.415 91.860 43.605 ;
        RECT 96.290 43.415 96.460 43.605 ;
        RECT 102.725 43.435 102.895 43.605 ;
        RECT 105.025 43.455 105.195 43.605 ;
        RECT 105.945 43.435 106.115 43.605 ;
        RECT 107.325 43.415 107.495 43.605 ;
        RECT 110.545 43.415 110.715 43.605 ;
        RECT 112.845 43.415 113.015 43.605 ;
        RECT 114.230 43.415 114.400 43.605 ;
        RECT 118.365 43.415 118.535 43.605 ;
        RECT 123.895 43.460 124.055 43.570 ;
      LAYER nwell ;
        RECT -0.190 42.165 97.135 42.215 ;
        RECT 98.760 42.165 124.850 42.215 ;
        RECT -0.190 39.435 124.850 42.165 ;
        RECT -0.190 39.385 96.675 39.435 ;
        RECT 98.300 39.385 124.850 39.435 ;
        RECT -0.190 36.725 97.135 36.775 ;
        RECT 98.760 36.725 124.850 36.775 ;
        RECT -0.190 33.995 124.850 36.725 ;
        RECT -0.190 33.945 96.675 33.995 ;
        RECT 98.300 33.945 124.850 33.995 ;
        RECT -0.190 31.285 97.135 31.335 ;
        RECT 98.760 31.285 124.850 31.335 ;
        RECT -0.190 28.555 124.850 31.285 ;
        RECT -0.190 28.505 96.675 28.555 ;
        RECT 98.300 28.505 124.850 28.555 ;
        RECT -0.190 25.845 97.135 25.895 ;
        RECT 98.760 25.845 124.850 25.895 ;
        RECT -0.190 23.115 124.850 25.845 ;
        RECT -0.190 23.065 96.675 23.115 ;
        RECT 98.300 23.065 124.850 23.115 ;
        RECT -0.190 20.405 97.135 20.455 ;
        RECT 98.760 20.405 124.850 20.455 ;
        RECT -0.190 17.675 124.850 20.405 ;
        RECT -0.190 17.625 96.675 17.675 ;
        RECT 98.300 17.625 124.850 17.675 ;
        RECT -0.190 14.965 97.135 15.015 ;
        RECT 98.760 14.965 124.850 15.015 ;
        RECT -0.190 12.235 124.850 14.965 ;
        RECT -0.190 12.185 96.675 12.235 ;
        RECT 98.300 12.185 124.850 12.235 ;
        RECT -0.190 9.525 97.135 9.575 ;
        RECT 98.760 9.525 124.850 9.575 ;
        RECT -0.190 6.795 124.850 9.525 ;
        RECT -0.190 6.745 96.675 6.795 ;
        RECT 98.300 6.745 124.850 6.795 ;
        RECT -0.190 4.085 97.135 4.135 ;
        RECT 98.760 4.085 124.850 4.135 ;
        RECT -0.190 1.355 124.850 4.085 ;
        RECT -0.190 1.305 96.675 1.355 ;
        RECT 98.300 1.305 124.850 1.355 ;
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 7.510 -0.085 7.680 0.105 ;
        RECT 12.105 -0.085 12.275 0.105 ;
        RECT 19.470 -0.085 19.640 0.105 ;
        RECT 24.065 -0.085 24.235 0.105 ;
        RECT 31.430 -0.085 31.600 0.105 ;
        RECT 36.025 -0.085 36.195 0.105 ;
        RECT 43.390 -0.085 43.560 0.105 ;
        RECT 47.985 -0.085 48.155 0.105 ;
        RECT 55.350 -0.085 55.520 0.105 ;
        RECT 59.945 -0.085 60.115 0.105 ;
        RECT 67.310 -0.085 67.480 0.105 ;
        RECT 71.905 -0.085 72.075 0.105 ;
        RECT 79.270 -0.085 79.440 0.105 ;
        RECT 83.865 -0.085 84.035 0.105 ;
        RECT 91.230 -0.085 91.400 0.105 ;
        RECT 95.830 -0.085 96.000 0.105 ;
        RECT 102.265 -0.085 102.435 0.085 ;
        RECT 104.565 -0.085 104.735 0.065 ;
        RECT 105.485 -0.085 105.655 0.085 ;
        RECT 106.865 -0.085 107.035 0.105 ;
        RECT 110.085 -0.085 110.255 0.105 ;
        RECT 112.385 -0.085 112.555 0.105 ;
        RECT 114.225 -0.085 114.395 0.105 ;
        RECT 119.745 -0.085 119.915 0.105 ;
        RECT 121.590 -0.085 121.760 0.105 ;
      LAYER li1 ;
        RECT 0.000 43.435 124.660 43.605 ;
      LAYER li1 ;
        RECT 0.000 0.085 124.660 43.435 ;
      LAYER li1 ;
        RECT 0.000 -0.085 124.660 0.085 ;
      LAYER met1 ;
        RECT 0.145 43.435 124.515 43.760 ;
        RECT 0.425 43.000 124.235 43.435 ;
        RECT 0.085 41.320 124.515 43.000 ;
        RECT 0.425 40.280 124.235 41.320 ;
        RECT 0.085 38.600 124.515 40.280 ;
        RECT 0.425 37.560 124.235 38.600 ;
        RECT 0.085 35.880 124.515 37.560 ;
        RECT 0.425 34.840 124.235 35.880 ;
        RECT 0.085 33.160 124.515 34.840 ;
        RECT 0.425 32.120 124.235 33.160 ;
        RECT 0.085 30.440 124.515 32.120 ;
        RECT 0.425 29.400 124.235 30.440 ;
        RECT 0.085 27.720 124.515 29.400 ;
        RECT 0.425 26.680 124.235 27.720 ;
        RECT 0.085 25.000 124.515 26.680 ;
        RECT 0.425 23.960 124.235 25.000 ;
        RECT 0.085 22.280 124.515 23.960 ;
        RECT 0.425 21.240 124.235 22.280 ;
        RECT 0.085 19.560 124.515 21.240 ;
        RECT 0.425 18.520 124.235 19.560 ;
        RECT 0.085 16.840 124.515 18.520 ;
        RECT 0.425 15.800 124.235 16.840 ;
        RECT 0.085 14.120 124.515 15.800 ;
        RECT 0.425 13.080 124.235 14.120 ;
        RECT 0.085 11.400 124.515 13.080 ;
        RECT 0.425 10.360 124.235 11.400 ;
        RECT 0.085 8.680 124.515 10.360 ;
        RECT 0.425 7.640 124.235 8.680 ;
        RECT 0.085 5.960 124.515 7.640 ;
        RECT 0.425 4.920 124.235 5.960 ;
        RECT 0.085 3.240 124.515 4.920 ;
        RECT 0.425 2.200 124.235 3.240 ;
        RECT 0.085 0.520 124.515 2.200 ;
        RECT 0.425 0.085 124.235 0.520 ;
        RECT 0.145 -0.240 124.515 0.085 ;
      LAYER met2 ;
        RECT 41.150 43.520 42.690 43.705 ;
        RECT 92.350 43.520 93.890 43.705 ;
        RECT 1.940 41.240 6.710 43.520 ;
        RECT 7.550 41.240 14.070 43.520 ;
        RECT 14.910 41.240 21.430 43.520 ;
        RECT 22.270 41.240 28.790 43.520 ;
        RECT 29.630 41.240 36.150 43.520 ;
        RECT 36.990 41.240 43.510 43.520 ;
        RECT 44.350 41.240 50.870 43.520 ;
        RECT 51.710 41.240 58.230 43.520 ;
        RECT 59.070 41.240 65.590 43.520 ;
        RECT 66.430 41.240 72.950 43.520 ;
        RECT 73.790 41.240 80.310 43.520 ;
        RECT 81.150 41.240 87.670 43.520 ;
        RECT 88.510 41.240 95.030 43.520 ;
        RECT 95.870 41.240 102.390 43.520 ;
        RECT 103.230 41.240 109.750 43.520 ;
        RECT 110.590 41.240 117.110 43.520 ;
        RECT 117.950 41.240 124.100 43.520 ;
        RECT 1.940 0.000 124.100 41.240 ;
        RECT 41.150 -0.185 42.690 0.000 ;
        RECT 92.350 -0.185 93.890 0.000 ;
      LAYER met3 ;
        RECT 41.130 43.520 42.710 43.685 ;
        RECT 92.330 43.520 93.910 43.685 ;
        RECT 11.105 37.760 122.660 43.520 ;
        RECT 11.105 36.360 122.260 37.760 ;
        RECT 11.105 32.320 122.660 36.360 ;
        RECT 11.105 30.920 122.260 32.320 ;
        RECT 11.105 26.880 122.660 30.920 ;
        RECT 11.105 25.480 122.260 26.880 ;
        RECT 11.105 21.440 122.660 25.480 ;
        RECT 11.105 20.040 122.260 21.440 ;
        RECT 11.105 16.000 122.660 20.040 ;
        RECT 11.105 14.600 122.260 16.000 ;
        RECT 11.105 10.560 122.660 14.600 ;
        RECT 11.105 9.160 122.260 10.560 ;
        RECT 11.105 5.120 122.660 9.160 ;
        RECT 11.105 3.720 122.260 5.120 ;
        RECT 11.105 0.000 122.660 3.720 ;
        RECT 41.130 -0.165 42.710 0.000 ;
        RECT 92.330 -0.165 93.910 0.000 ;
  END
END RAM16
END LIBRARY

